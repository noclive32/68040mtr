--==========================> Motorola 68040 <===========================--
-- RESET_IRQ_HANDLER.VHD	
-- Engineer:	Kevin Phillipson
-- Date:		10/28/2007									Revision:10.28.07
-- Description: Generates interrupt condition signal and correct interrupt
-- vector.  It also immplements the reset logic
--
-- 
-- These signals cause a system reset and are nonmaskable. The interrupt
-- vectors are implemented here. A list of the signals and vectors is
-- provided below:
--
--		nreset			FFFE	reset
--		clm_sig			FFFC	clock monitor timeout
--		cop_sig			FFFA	cop timeout
--
-- These interrupt vectors are generated by opcodes and are therefore
-- hardcoded into the microcode and are not implemented here:
--
--		invalid opcode	FFF8	illegal opcode trap
--		opcode 0x3F		FFF6	swi
--
-- These interrupt vectors are implemented here. They are maskable by the
-- X and I bits in the CCR. A list of the signals and vectors is provided
-- below:
--
--		dev_irq( 0)		FFF4	xirq pin (pseudo non-maskable interrupt)
--		dev_irq( 1)		FFF2	irq (external pin or parallel i/o)
--		dev_irq( 2)		FFF0	real time interrupt
--		dev_irq( 3)		FFEE	timer input capture 1
--		dev_irq( 4)		FFEC	timer input capture 2
--		dev_irq( 5)		FFEA	timer input capture 3
--		dev_irq( 6)		FFE8	timer output compare 1
--		dev_irq( 7)		FFE6	timer output compare 2
--		dev_irq( 8)		FFE4	timer output compare 3
--		dev_irq( 9)		FFE2	timer output compare 4
--		dev_irq(10)		FFE0	timer output compare 5
--		dev_irq(11)		FFDE	timer overflow
--		dev_irq(12)		FFDC	pulse accumulator overflow
--		dev_irq(13)		FFDA	pulse accumulator input edge
--		dev_irq(14)		FFD8	SPI serial transfer complete
--		dev_irq(15)		FFD6	SCI serial system
-- 
--==========================================================================--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity reset_irq_handler is

--============================> Port Map <==================================--

port
(
	----------------------------------------> Inputs
	--
	nreset		:	in	std_logic;	-- Negative Logic System Reset

	clk			:	in	std_logic;	-- System Clock
	
	cop_sig		:	in	std_logic;	-- Computer Operating Properly Reset Signal
	clm_sig		:	in	std_logic;	-- Clock Monitor Reset Signal

	ipsel		:	in	std_logic_vector( 3 downto  0);	-- Interrupt Priority Select

	ccr_data	:	in	std_logic_vector( 7 downto  0);	-- Condition Code Register Flags
	
	dev_irq		:	in	std_logic_vector(15 downto  0); -- Device Interrupt ReQuests
	--
	---------------------------------------->


	----------------------------------------> Outputs
	--
	sys_rst		:	out	std_logic;

	stop_cond	:	out	std_logic;

	irq_cond	:	out	std_logic;

	set_x_msk	:	out	std_logic;
	
	irq_vec		:	out	std_logic_vector(15 downto  0)
	--
	----------------------------------------< 

);

--==========================================================================--

end reset_irq_handler;

architecture behavior of reset_irq_handler is 

--==============================> Signals <=================================--


constant	RST_VEC			:	std_logic_vector( 7 downto  0)	:=	x"FE";	-- clock monitor timeout
constant	CLM_VEC			:	std_logic_vector( 7 downto  0)	:=	x"FC";	-- clock monitor timeout
constant	COP_VEC			:	std_logic_vector( 7 downto  0)	:=	x"FA";	-- cop timeout
constant	DEV_00_VEC		:	std_logic_vector( 7 downto  0)	:=	x"F4";	-- xirq pin (pseudo non-maskable interrupt)
constant	DEV_01_VEC		:	std_logic_vector( 7 downto  0)	:=	x"F2";	-- irq (external pin or parallel i/o)
constant	DEV_02_VEC		:	std_logic_vector( 7 downto  0)	:=	x"F0";	-- real time interrupt
constant	DEV_03_VEC		:	std_logic_vector( 7 downto  0)	:=	x"EE";	-- timer input capture 1
constant	DEV_04_VEC		:	std_logic_vector( 7 downto  0)	:=	x"EC";	-- timer input capture 2
constant	DEV_05_VEC		:	std_logic_vector( 7 downto  0)	:=	x"EA";	-- timer input capture 3
constant	DEV_06_VEC		:	std_logic_vector( 7 downto  0)	:=	x"E8";	-- timer output compare 1
constant	DEV_07_VEC		:	std_logic_vector( 7 downto  0)	:=	x"E6";	-- timer output compare 2
constant	DEV_08_VEC		:	std_logic_vector( 7 downto  0)	:=	x"E4";	-- timer output compare 3
constant	DEV_09_VEC		:	std_logic_vector( 7 downto  0)	:=	x"E2";	-- timer output compare 4
constant	DEV_10_VEC		:	std_logic_vector( 7 downto  0)	:=	x"E0";	-- timer output compare 5
constant	DEV_11_VEC		:	std_logic_vector( 7 downto  0)	:=	x"DE";	-- timer overflow
constant	DEV_12_VEC		:	std_logic_vector( 7 downto  0)	:=	x"DC";	-- pulse accumulator overflow
constant	DEV_13_VEC		:	std_logic_vector( 7 downto  0)	:=	x"DA";	-- pulse accumulator input edge
constant	DEV_14_VEC		:	std_logic_vector( 7 downto  0)	:=	x"D8";	-- SPI serial transfer complete
constant	DEV_15_VEC		:	std_logic_vector( 7 downto  0)	:=	x"D6";	-- SCI serial system

signal		ccr_x			:	std_logic;
signal		ccr_i			:	std_logic;
signal		ccr_s			:	std_logic;

signal		set_x_msk_nxt	:	std_logic;
signal		set_x_msk_reg	:	std_logic;

signal		irq_cond_nxt	:	std_logic;
signal		irq_cond_reg	:	std_logic;

signal		stop_cond_reg	:	std_logic;

signal		irq_vec_nxt		:	std_logic_vector( 7 downto  0);
signal		irq_vec_reg		:	std_logic_vector( 7 downto  0);

signal		priority_irq	:	std_logic;
signal		priority_vec	:	std_logic_vector( 7 downto  0);

signal		sys_rst_reg		:	std_logic;
signal		rst_reg			:	std_logic;
signal		clm_reg			:	std_logic;
signal		cop_reg			:	std_logic;
signal		rst_sreg		:	std_logic_vector( 1 downto  0);


--==========================================================================--

begin

--===========================> Architecture <===============================--


----------------------------------------> Reset Logic
--

process
(
	clk,
	nreset,
	clm_sig,
	cop_sig,
	rst_sreg
)
begin

	if (clk'event and clk = '1') then
	
		--2bit shift reg
		rst_sreg(0)	<= not nreset;
		rst_sreg(1)	<= rst_sreg(0);

		--Synchronized System Reset for internal and external devices
		if (rst_sreg = "11" or clm_sig = '1' or cop_sig = '1') then
			sys_rst_reg	<=	'1';
		else
			sys_rst_reg	<=	'0';
		end if;

		--Synchronized External Reset for interrupt vector logic
		if (rst_sreg = "11") then
			rst_reg	<= '1';
		else
			rst_reg	<= '0';
		end if;
	
		--Synchronized COP & CLM for interrupt vector logic
		cop_reg	<=	cop_sig;
		clm_reg	<=	clm_sig;
	
	end if;

end process;

sys_rst	<=	sys_rst_reg;
--
----------------------------------------<


----------------------------------------> Stop Instruction Condition Logic
--

ccr_s	<=	ccr_data(7);

process
(
	clk,
	ccr_i,
	ccr_s,
	dev_irq
)
begin

	if (clk'event and clk = '1') then

		-- if (ccr_s=1 or xirq=1 or (ccr_i=0 and irq=1))
		if (ccr_s='1' or dev_irq(0)='1' or (ccr_i='1' and dev_irq(1)='1')) then
			-- don't stop
			stop_cond_reg	<=	'0';
		else
			-- stop
			stop_cond_reg	<=	'1';
		end if;
	
	end if;

end process;

stop_cond	<=	stop_cond_reg;
--
----------------------------------------<

----------------------------------------> Interrupt Decoding Logic
--

ccr_i	<=	ccr_data(4);
ccr_x	<=	ccr_data(6);

with ipsel select
priority_irq	<=
	dev_irq(11)	when x"0",	-- timer overflow
	dev_irq(12)	when x"1",	-- pulse accumulator overflow
	dev_irq(13)	when x"2",	-- pulse accumulator input edge
	dev_irq(14)	when x"3",	-- SPI serial transfer complete
	dev_irq(15)	when x"4",	-- SCI serial system
	dev_irq( 1)	when x"5",	-- reserved (default to irq)
	dev_irq( 1)	when x"6",	-- irq (external pin or parallel i/o)
	dev_irq( 2)	when x"7",	-- real time interrupt
	dev_irq( 3)	when x"8",	-- timer input capture 1
	dev_irq( 4)	when x"9",	-- timer input capture 2
	dev_irq( 5)	when x"A",	-- timer input capture 3
	dev_irq( 6)	when x"B",	-- timer output compare 1
	dev_irq( 7)	when x"C",	-- timer output compare 2
	dev_irq( 8)	when x"D",	-- timer output compare 3
	dev_irq( 9)	when x"E",	-- timer output compare 4
	dev_irq(10)	when others; --x"F" timer output compare 5

with ipsel select
priority_vec	<=
	DEV_11_VEC	when x"0",	-- timer overflow
	DEV_12_VEC	when x"1",	-- pulse accumulator overflow
	DEV_13_VEC	when x"2",	-- pulse accumulator input edge
	DEV_14_VEC	when x"3",	-- SPI serial transfer complete
	DEV_15_VEC	when x"4",	-- SCI serial system
	DEV_01_VEC	when x"5",	-- reserved (default to irq)
	DEV_01_VEC	when x"6",	-- irq (external pin or parallel i/o)
	DEV_02_VEC	when x"7",	-- real time interrupt
	DEV_03_VEC	when x"8",	-- timer input capture 1
	DEV_04_VEC	when x"9",	-- timer input capture 2
	DEV_05_VEC	when x"A",	-- timer input capture 3
	DEV_06_VEC	when x"B",	-- timer output compare 1
	DEV_07_VEC	when x"C",	-- timer output compare 2
	DEV_08_VEC	when x"D",	-- timer output compare 3
	DEV_09_VEC	when x"E",	-- timer output compare 4
	DEV_10_VEC	when others; --x"F" timer output compare 5

process
(
	rst_reg,
	cop_reg,
	clm_reg,
	set_x_msk_reg,
	irq_vec_reg,
	ccr_i,
	ccr_x,
	priority_vec,
	priority_irq,
	dev_irq
)
begin

	-- Default next values if no interrupt
	irq_cond_nxt	<=	'0';
	set_x_msk_nxt	<=	set_x_msk_reg;
	irq_vec_nxt		<=	irq_vec_reg;

	if (rst_reg = '1') then	-- External Reset
		irq_cond_nxt	<=	'0';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	RST_VEC;

	elsif (clm_reg = '1') then	-- Clock Monitor Reset
		irq_cond_nxt	<=	'0';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	CLM_VEC;
	
	elsif (cop_reg = '1') then	-- Computer Operating Properly Reset
		irq_cond_nxt	<=	'0';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	COP_VEC;

	elsif (dev_irq( 0) = '1' and ccr_x = '0') then -- xirq pin (pseudo non-maskable interrupt)
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'1';
		irq_vec_nxt		<=	DEV_00_VEC;

	elsif (priority_irq = '1' and ccr_i = '0') then	-- priority irq (selected by ipsel)
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	priority_vec;

	elsif (dev_irq( 1) = '1' and ccr_i = '0') then	-- irq (external pin or parallel i/o)
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_01_VEC;

	elsif (dev_irq( 2) = '1' and ccr_i = '0') then	-- real time interrupt
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_02_VEC;
	
	elsif (dev_irq( 3) = '1' and ccr_i = '0') then	-- timer input capture 1
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_03_VEC;
	
	elsif (dev_irq( 4) = '1' and ccr_i = '0') then	-- timer input capture 2
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_04_VEC;
	
	elsif (dev_irq( 5) = '1' and ccr_i = '0') then	-- timer input capture 3
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_05_VEC;
	
	elsif (dev_irq( 6) = '1' and ccr_i = '0') then	-- timer output compare 1
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_06_VEC;

	elsif (dev_irq( 7) = '1' and ccr_i = '0') then	-- timer output compare 2
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_07_VEC;

	elsif (dev_irq( 8) = '1' and ccr_i = '0') then	-- timer output compare 3
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_08_VEC;
	
	elsif (dev_irq( 9) = '1' and ccr_i = '0') then	-- timer output compare 4
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_09_VEC;
	
	elsif (dev_irq(10) = '1' and ccr_i = '0') then	-- timer output compare 5
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_10_VEC;
	
	elsif (dev_irq(11) = '1' and ccr_i = '0') then	-- timer overflow
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_11_VEC;
	
	elsif (dev_irq(12) = '1' and ccr_i = '0') then	-- pulse accumulator overflow
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_12_VEC;
	
	elsif (dev_irq(13) = '1' and ccr_i = '0') then	-- pulse accumulator input edge
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_13_VEC;
	
	elsif (dev_irq(14) = '1' and ccr_i = '0') then	-- SPI serial transfer complete
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_14_VEC;
	
	elsif (dev_irq(15) = '1' and ccr_i = '0') then	-- SCI serial system
		irq_cond_nxt	<=	'1';
		set_x_msk_nxt	<=	'0';
		irq_vec_nxt		<=	DEV_15_VEC;
	end if;

end process;

process
(
	clk,
	irq_cond_nxt,
	set_x_msk_nxt,
	irq_vec_nxt
)
begin

	if (clk'event and clk = '1') then
	
		irq_cond_reg	<=	irq_cond_nxt;
		set_x_msk_reg	<=	set_x_msk_nxt;
		irq_vec_reg		<=	irq_vec_nxt;

	end if;

end process;

set_x_msk	<=	set_x_msk_reg;
irq_cond	<=	irq_cond_reg;
irq_vec		<=	x"FF" & irq_vec_reg;
--
----------------------------------------<


--==========================================================================--
end behavior;






